LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;

entity game_lx_ram is
port(
	reset : in std_logic;
	died : out std_logic;
	clock_s : in std_logic;
	print : inout std_logic;
	clk : in std_logic;
	size : in integer range 40 downto 4;
	applexout : in integer range 63 downto 0;
	appleyout : in integer range 31 downto 0;
	xout : in integer range 63 downto 0;
	yout : in integer range 31 downto 0;
	lineout : out std_logic_vector(127 downto 0)
);
end game_lx_ram;

architecture game_lx_ram_ar of game_lx_ram is
signal en : integer range 41 downto 0;
begin
process(clk,clock_s)
variable xtemp : integer range 63 downto 0;
variable	ytemp : integer range 31 downto 0;
variable delay : integer range 4 downto 0;
variable num : integer range 16 downto 0;
variable linenum : integer range 63 downto 0;
variable l0,l1,l2,l3,l4,l5,l6,l7,l8,l9,l10,l11,l12,l13,l14,l15,l16,l17,l18,l19,l20,l21,l22,l23,l24,l25,l26,l27,l28,l29,l30,l31,l32,l33,l34,l35,l36,l37,l38,l39,l40,l41,l42,l43,l44,l45,l46,l47,l48,l49,l50,l51,l52,l53,l54,l55,l56,l57,l58,l59,l60,l61,l62,l63 : std_logic_vector(0 to 127);
begin
if(clock_s='0')then
en<=size+1;
if(reset='1')then
print<='0';
died<='0';
end if;
	delay:=3;
	linenum:=0;
	num:=16;
l0:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l1:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l2:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l3:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l4:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l5:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l6:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l7:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l8:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l9:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l10:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l11:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l12:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l13:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l14:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l15:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l16:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l17:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l18:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l19:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l20:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l21:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l22:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l23:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l24:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l25:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l26:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l27:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l28:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l29:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l30:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l31:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l32:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l33:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l34:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l35:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l36:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l37:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l38:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l39:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l40:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l41:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l42:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l43:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l44:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l45:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l46:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l47:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l48:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l49:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l50:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l51:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l52:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l53:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l54:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l55:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l56:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l57:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l58:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l59:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l60:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l61:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l62:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
l63:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
elsif(clock_s='1')then 
	if(clk'event and clk='1')then
		if en>1 then
		
		ytemp:=yout;
		xtemp:=xout;
		elsif en=1 then
		ytemp:=appleyout;
		xtemp:=applexout;
		
		end if;
		if(en>0)then
		en<=en-1;
	case ytemp is
	when 0 =>
if l0(2*xtemp)='1' then
died<='1';
end if;
l0(2*xtemp):='1';
l0(2*xtemp+1):='1';
l1(2*xtemp):='1';
l1(2*xtemp+1):='1';
when 1 =>
if l2(2*xtemp)='1' then
died<='1';
end if;
l2(2*xtemp):='1';
l2(2*xtemp+1):='1';
l3(2*xtemp):='1';
l3(2*xtemp+1):='1';
when 2 =>
if l4(2*xtemp)='1' then
died<='1';
end if;
l4(2*xtemp):='1';
l4(2*xtemp+1):='1';
l5(2*xtemp):='1';
l5(2*xtemp+1):='1';
when 3 =>
if l6(2*xtemp)='1' then
died<='1';
end if;
l6(2*xtemp):='1';
l6(2*xtemp+1):='1';
l7(2*xtemp):='1';
l7(2*xtemp+1):='1';
when 4 =>
if l8(2*xtemp)='1' then
died<='1';
end if;
l8(2*xtemp):='1';
l8(2*xtemp+1):='1';
l9(2*xtemp):='1';
l9(2*xtemp+1):='1';
when 5 =>
if l10(2*xtemp)='1' then
died<='1';
end if;
l10(2*xtemp):='1';
l10(2*xtemp+1):='1';
l11(2*xtemp):='1';
l11(2*xtemp+1):='1';
when 6 =>
if l12(2*xtemp)='1' then
died<='1';
end if;
l12(2*xtemp):='1';
l12(2*xtemp+1):='1';
l13(2*xtemp):='1';
l13(2*xtemp+1):='1';
when 7 =>
if l14(2*xtemp)='1' then
died<='1';
end if;
l14(2*xtemp):='1';
l14(2*xtemp+1):='1';
l15(2*xtemp):='1';
l15(2*xtemp+1):='1';
when 8 =>
if l16(2*xtemp)='1' then
died<='1';
end if;
l16(2*xtemp):='1';
l16(2*xtemp+1):='1';
l17(2*xtemp):='1';
l17(2*xtemp+1):='1';
when 9 =>
if l18(2*xtemp)='1' then
died<='1';
end if;
l18(2*xtemp):='1';
l18(2*xtemp+1):='1';
l19(2*xtemp):='1';
l19(2*xtemp+1):='1';
when 10 =>
if l20(2*xtemp)='1' then
died<='1';
end if;
l20(2*xtemp):='1';
l20(2*xtemp+1):='1';
l21(2*xtemp):='1';
l21(2*xtemp+1):='1';
when 11 =>
if l22(2*xtemp)='1' then
died<='1';
end if;
l22(2*xtemp):='1';
l22(2*xtemp+1):='1';
l23(2*xtemp):='1';
l23(2*xtemp+1):='1';
when 12 =>
if l24(2*xtemp)='1' then
died<='1';
end if;
l24(2*xtemp):='1';
l24(2*xtemp+1):='1';
l25(2*xtemp):='1';
l25(2*xtemp+1):='1';
when 13 =>
if l26(2*xtemp)='1' then
died<='1';
end if;
l26(2*xtemp):='1';
l26(2*xtemp+1):='1';
l27(2*xtemp):='1';
l27(2*xtemp+1):='1';
when 14 =>
if l28(2*xtemp)='1' then
died<='1';
end if;
l28(2*xtemp):='1';
l28(2*xtemp+1):='1';
l29(2*xtemp):='1';
l29(2*xtemp+1):='1';
when 15 =>
if l30(2*xtemp)='1' then
died<='1';
end if;
l30(2*xtemp):='1';
l30(2*xtemp+1):='1';
l31(2*xtemp):='1';
l31(2*xtemp+1):='1';
when 16 =>
if l32(2*xtemp)='1' then
died<='1';
end if;
l32(2*xtemp):='1';
l32(2*xtemp+1):='1';
l33(2*xtemp):='1';
l33(2*xtemp+1):='1';
when 17 =>
if l34(2*xtemp)='1' then
died<='1';
end if;
l34(2*xtemp):='1';
l34(2*xtemp+1):='1';
l35(2*xtemp):='1';
l35(2*xtemp+1):='1';
when 18 =>
if l36(2*xtemp)='1' then
died<='1';
end if;
l36(2*xtemp):='1';
l36(2*xtemp+1):='1';
l37(2*xtemp):='1';
l37(2*xtemp+1):='1';
when 19 =>
if l38(2*xtemp)='1' then
died<='1';
end if;
l38(2*xtemp):='1';
l38(2*xtemp+1):='1';
l39(2*xtemp):='1';
l39(2*xtemp+1):='1';
when 20 =>
if l40(2*xtemp)='1' then
died<='1';
end if;
l40(2*xtemp):='1';
l40(2*xtemp+1):='1';
l41(2*xtemp):='1';
l41(2*xtemp+1):='1';
when 21 =>
if l42(2*xtemp)='1' then
died<='1';
end if;
l42(2*xtemp):='1';
l42(2*xtemp+1):='1';
l43(2*xtemp):='1';
l43(2*xtemp+1):='1';
when 22 =>
if l44(2*xtemp)='1' then
died<='1';
end if;
l44(2*xtemp):='1';
l44(2*xtemp+1):='1';
l45(2*xtemp):='1';
l45(2*xtemp+1):='1';
when 23 =>
if l46(2*xtemp)='1' then
died<='1';
end if;
l46(2*xtemp):='1';
l46(2*xtemp+1):='1';
l47(2*xtemp):='1';
l47(2*xtemp+1):='1';
when 24 =>
if l48(2*xtemp)='1' then
died<='1';
end if;
l48(2*xtemp):='1';
l48(2*xtemp+1):='1';
l49(2*xtemp):='1';
l49(2*xtemp+1):='1';
when 25 =>
if l50(2*xtemp)='1' then
died<='1';
end if;
l50(2*xtemp):='1';
l50(2*xtemp+1):='1';
l51(2*xtemp):='1';
l51(2*xtemp+1):='1';
when 26 =>
if l52(2*xtemp)='1' then
died<='1';
end if;
l52(2*xtemp):='1';
l52(2*xtemp+1):='1';
l53(2*xtemp):='1';
l53(2*xtemp+1):='1';
when 27 =>
if l54(2*xtemp)='1' then
died<='1';
end if;
l54(2*xtemp):='1';
l54(2*xtemp+1):='1';
l55(2*xtemp):='1';
l55(2*xtemp+1):='1';
when 28 =>
if l56(2*xtemp)='1' then
died<='1';
end if;
l56(2*xtemp):='1';
l56(2*xtemp+1):='1';
l57(2*xtemp):='1';
l57(2*xtemp+1):='1';
when 29 =>
if l58(2*xtemp)='1' then
died<='1';
end if;
l58(2*xtemp):='1';
l58(2*xtemp+1):='1';
l59(2*xtemp):='1';
l59(2*xtemp+1):='1';
when 30 =>
if l60(2*xtemp)='1' then
died<='1';
end if;
l60(2*xtemp):='1';
l60(2*xtemp+1):='1';
l61(2*xtemp):='1';
l61(2*xtemp+1):='1';
when 31 =>
if l62(2*xtemp)='1' then
died<='1';
end if;
l62(2*xtemp):='1';
l62(2*xtemp+1):='1';
l63(2*xtemp):='1';
l63(2*xtemp+1):='1';


	end case;
		end if;
		if(en=0)then 
		print<='1';
		end if;
		
		if(print='1')then
		if delay>0 then 
		delay:=delay-1;
		elsif num=16 then
		num:=0;
		
			case linenum is
			when 0=>
lineout<=l0;
when 1=>
lineout<=l1;
when 2=>
lineout<=l2;
when 3=>
lineout<=l3;
when 4=>
lineout<=l4;
when 5=>
lineout<=l5;
when 6=>
lineout<=l6;
when 7=>
lineout<=l7;
when 8=>
lineout<=l8;
when 9=>
lineout<=l9;
when 10=>
lineout<=l10;
when 11=>
lineout<=l11;
when 12=>
lineout<=l12;
when 13=>
lineout<=l13;
when 14=>
lineout<=l14;
when 15=>
lineout<=l15;
when 16=>
lineout<=l16;
when 17=>
lineout<=l17;
when 18=>
lineout<=l18;
when 19=>
lineout<=l19;
when 20=>
lineout<=l20;
when 21=>
lineout<=l21;
when 22=>
lineout<=l22;
when 23=>
lineout<=l23;
when 24=>
lineout<=l24;
when 25=>
lineout<=l25;
when 26=>
lineout<=l26;
when 27=>
lineout<=l27;
when 28=>
lineout<=l28;
when 29=>
lineout<=l29;
when 30=>
lineout<=l30;
when 31=>
lineout<=l31;
when 32=>
lineout<=l32;
when 33=>
lineout<=l33;
when 34=>
lineout<=l34;
when 35=>
lineout<=l35;
when 36=>
lineout<=l36;
when 37=>
lineout<=l37;
when 38=>
lineout<=l38;
when 39=>
lineout<=l39;
when 40=>
lineout<=l40;
when 41=>
lineout<=l41;
when 42=>
lineout<=l42;
when 43=>
lineout<=l43;
when 44=>
lineout<=l44;
when 45=>
lineout<=l45;
when 46=>
lineout<=l46;
when 47=>
lineout<=l47;
when 48=>
lineout<=l48;
when 49=>
lineout<=l49;
when 50=>
lineout<=l50;
when 51=>
lineout<=l51;
when 52=>
lineout<=l52;
when 53=>
lineout<=l53;
when 54=>
lineout<=l54;
when 55=>
lineout<=l55;
when 56=>
lineout<=l56;
when 57=>
lineout<=l57;
when 58=>
lineout<=l58;
when 59=>
lineout<=l59;
when 60=>
lineout<=l60;
when 61=>
lineout<=l61;
when 62=>
lineout<=l62;
when 63=>
lineout<=l63;
			end case;
		if linenum<64 then
			linenum:=linenum+1;
		else print<='0';
		end if;
		
		elsif num<16 then
			num:=num+1;
			
		end if;
		end if;
	end if;	
	end if;
end process;
end game_lx_ram_ar;